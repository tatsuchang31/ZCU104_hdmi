library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package type_pack is

constant RAM_DATALENGTH	: INTEGER := 48;
constant RAM_ADDRESS	: INTEGER := 16384;
constant RAM_ADDRESSBIT	: INTEGER := 14;

constant H_POS	: INTEGER := 1920;
constant V_POS	: INTEGER := 1080;

end package type_pack;